--Command Processor 
--Daryl White and Alexander Hamilton

--code goes here